library ieee;
use ieee.std_logic_1164.all;

entity neander is
    port(
        cl, clk : in std_logic;
    );
end entity;

architecture cha_mate of neander is
    component ula is
        port(

        );
    end component;

    component memory is
        port(

        );
    end component;
begin

end architecture;