entity uc_control is
    --port(

    --);
end entity;

architecture hohoho_o_cacetinho of uc_control is

begin

end architecture;