entity decoder is
    port(

    );
end entity;



architecture minipizzas of decoder is

begin

end architecture;