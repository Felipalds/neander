entity pc is
    port(

    );
end entity;

architecture brigadeiros of pc is

begin

end architecture;